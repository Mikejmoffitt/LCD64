library ieee;
use ieee.std_logic_1164.all;

entity gamma_curver is
port (
	sig_in: in std_logic_vector(7 downto 0);
	sig_out: out std_logic_vector(7 downto 0));
end entity;

architecture behavioral of gamma_curver is
begin
	lookup: process(sig_in)
	begin
	if (sig_in = X"00") then
		sig_out <= X"00";
	elsif (sig_in = X"01") then
		sig_out <= X"00";
	elsif (sig_in = X"02") then
		sig_out <= X"01";
	elsif (sig_in = X"03") then
		sig_out <= X"01";
	elsif (sig_in = X"04") then
		sig_out <= X"02";
	elsif (sig_in = X"05") then
		sig_out <= X"02";
	elsif (sig_in = X"06") then
		sig_out <= X"03";
	elsif (sig_in = X"07") then
		sig_out <= X"03";
	elsif (sig_in = X"08") then
		sig_out <= X"04";
	elsif (sig_in = X"09") then
		sig_out <= X"04";
	elsif (sig_in = X"0A") then
		sig_out <= X"05";
	elsif (sig_in = X"0B") then
		sig_out <= X"05";
	elsif (sig_in = X"0C") then
		sig_out <= X"06";
	elsif (sig_in = X"0D") then
		sig_out <= X"06";
	elsif (sig_in = X"0E") then
		sig_out <= X"07";
	elsif (sig_in = X"0F") then
		sig_out <= X"07";
	elsif (sig_in = X"10") then
		sig_out <= X"08";
	elsif (sig_in = X"11") then
		sig_out <= X"08";
	elsif (sig_in = X"12") then
		sig_out <= X"09";
	elsif (sig_in = X"13") then
		sig_out <= X"09";
	elsif (sig_in = X"14") then
		sig_out <= X"0A";
	elsif (sig_in = X"15") then
		sig_out <= X"0A";
	elsif (sig_in = X"16") then
		sig_out <= X"0B";
	elsif (sig_in = X"17") then
		sig_out <= X"0B";
	elsif (sig_in = X"18") then
		sig_out <= X"0C";
	elsif (sig_in = X"19") then
		sig_out <= X"0C";
	elsif (sig_in = X"1A") then
		sig_out <= X"0D";
	elsif (sig_in = X"1B") then
		sig_out <= X"0D";
	elsif (sig_in = X"1C") then
		sig_out <= X"0E";
	elsif (sig_in = X"1D") then
		sig_out <= X"0F";
	elsif (sig_in = X"1E") then
		sig_out <= X"0F";
	elsif (sig_in = X"1F") then
		sig_out <= X"10";
	elsif (sig_in = X"20") then
		sig_out <= X"10";
	elsif (sig_in = X"21") then
		sig_out <= X"11";
	elsif (sig_in = X"22") then
		sig_out <= X"11";
	elsif (sig_in = X"23") then
		sig_out <= X"12";
	elsif (sig_in = X"24") then
		sig_out <= X"12";
	elsif (sig_in = X"25") then
		sig_out <= X"13";
	elsif (sig_in = X"26") then
		sig_out <= X"13";
	elsif (sig_in = X"27") then
		sig_out <= X"14";
	elsif (sig_in = X"28") then
		sig_out <= X"14";
	elsif (sig_in = X"29") then
		sig_out <= X"15";
	elsif (sig_in = X"2A") then
		sig_out <= X"16";
	elsif (sig_in = X"2B") then
		sig_out <= X"16";
	elsif (sig_in = X"2C") then
		sig_out <= X"17";
	elsif (sig_in = X"2D") then
		sig_out <= X"17";
	elsif (sig_in = X"2E") then
		sig_out <= X"18";
	elsif (sig_in = X"2F") then
		sig_out <= X"18";
	elsif (sig_in = X"30") then
		sig_out <= X"19";
	elsif (sig_in = X"31") then
		sig_out <= X"1A";
	elsif (sig_in = X"32") then
		sig_out <= X"1A";
	elsif (sig_in = X"33") then
		sig_out <= X"1B";
	elsif (sig_in = X"34") then
		sig_out <= X"1B";
	elsif (sig_in = X"35") then
		sig_out <= X"1C";
	elsif (sig_in = X"36") then
		sig_out <= X"1C";
	elsif (sig_in = X"37") then
		sig_out <= X"1D";
	elsif (sig_in = X"38") then
		sig_out <= X"1E";
	elsif (sig_in = X"39") then
		sig_out <= X"1E";
	elsif (sig_in = X"3A") then
		sig_out <= X"1F";
	elsif (sig_in = X"3B") then
		sig_out <= X"1F";
	elsif (sig_in = X"3C") then
		sig_out <= X"20";
	elsif (sig_in = X"3D") then
		sig_out <= X"21";
	elsif (sig_in = X"3E") then
		sig_out <= X"21";
	elsif (sig_in = X"3F") then
		sig_out <= X"22";
	elsif (sig_in = X"40") then
		sig_out <= X"22";
	elsif (sig_in = X"41") then
		sig_out <= X"23";
	elsif (sig_in = X"42") then
		sig_out <= X"24";
	elsif (sig_in = X"43") then
		sig_out <= X"24";
	elsif (sig_in = X"44") then
		sig_out <= X"25";
	elsif (sig_in = X"45") then
		sig_out <= X"26";
	elsif (sig_in = X"46") then
		sig_out <= X"26";
	elsif (sig_in = X"47") then
		sig_out <= X"27";
	elsif (sig_in = X"48") then
		sig_out <= X"27";
	elsif (sig_in = X"49") then
		sig_out <= X"28";
	elsif (sig_in = X"4A") then
		sig_out <= X"29";
	elsif (sig_in = X"4B") then
		sig_out <= X"29";
	elsif (sig_in = X"4C") then
		sig_out <= X"2A";
	elsif (sig_in = X"4D") then
		sig_out <= X"2B";
	elsif (sig_in = X"4E") then
		sig_out <= X"2B";
	elsif (sig_in = X"4F") then
		sig_out <= X"2C";
	elsif (sig_in = X"50") then
		sig_out <= X"2D";
	elsif (sig_in = X"51") then
		sig_out <= X"2D";
	elsif (sig_in = X"52") then
		sig_out <= X"2E";
	elsif (sig_in = X"53") then
		sig_out <= X"2F";
	elsif (sig_in = X"54") then
		sig_out <= X"2F";
	elsif (sig_in = X"55") then
		sig_out <= X"30";
	elsif (sig_in = X"56") then
		sig_out <= X"31";
	elsif (sig_in = X"57") then
		sig_out <= X"32";
	elsif (sig_in = X"58") then
		sig_out <= X"32";
	elsif (sig_in = X"59") then
		sig_out <= X"33";
	elsif (sig_in = X"5A") then
		sig_out <= X"34";
	elsif (sig_in = X"5B") then
		sig_out <= X"34";
	elsif (sig_in = X"5C") then
		sig_out <= X"35";
	elsif (sig_in = X"5D") then
		sig_out <= X"36";
	elsif (sig_in = X"5E") then
		sig_out <= X"37";
	elsif (sig_in = X"5F") then
		sig_out <= X"37";
	elsif (sig_in = X"60") then
		sig_out <= X"38";
	elsif (sig_in = X"61") then
		sig_out <= X"39";
	elsif (sig_in = X"62") then
		sig_out <= X"3A";
	elsif (sig_in = X"63") then
		sig_out <= X"3A";
	elsif (sig_in = X"64") then
		sig_out <= X"3B";
	elsif (sig_in = X"65") then
		sig_out <= X"3C";
	elsif (sig_in = X"66") then
		sig_out <= X"3D";
	elsif (sig_in = X"67") then
		sig_out <= X"3D";
	elsif (sig_in = X"68") then
		sig_out <= X"3E";
	elsif (sig_in = X"69") then
		sig_out <= X"3F";
	elsif (sig_in = X"6A") then
		sig_out <= X"40";
	elsif (sig_in = X"6B") then
		sig_out <= X"40";
	elsif (sig_in = X"6C") then
		sig_out <= X"41";
	elsif (sig_in = X"6D") then
		sig_out <= X"42";
	elsif (sig_in = X"6E") then
		sig_out <= X"43";
	elsif (sig_in = X"6F") then
		sig_out <= X"44";
	elsif (sig_in = X"70") then
		sig_out <= X"44";
	elsif (sig_in = X"71") then
		sig_out <= X"45";
	elsif (sig_in = X"72") then
		sig_out <= X"46";
	elsif (sig_in = X"73") then
		sig_out <= X"47";
	elsif (sig_in = X"74") then
		sig_out <= X"48";
	elsif (sig_in = X"75") then
		sig_out <= X"49";
	elsif (sig_in = X"76") then
		sig_out <= X"49";
	elsif (sig_in = X"77") then
		sig_out <= X"4A";
	elsif (sig_in = X"78") then
		sig_out <= X"4B";
	elsif (sig_in = X"79") then
		sig_out <= X"4C";
	elsif (sig_in = X"7A") then
		sig_out <= X"4D";
	elsif (sig_in = X"7B") then
		sig_out <= X"4E";
	elsif (sig_in = X"7C") then
		sig_out <= X"4F";
	elsif (sig_in = X"7D") then
		sig_out <= X"50";
	elsif (sig_in = X"7E") then
		sig_out <= X"50";
	elsif (sig_in = X"7F") then
		sig_out <= X"51";
	elsif (sig_in = X"80") then
		sig_out <= X"52";
	elsif (sig_in = X"81") then
		sig_out <= X"53";
	elsif (sig_in = X"82") then
		sig_out <= X"54";
	elsif (sig_in = X"83") then
		sig_out <= X"55";
	elsif (sig_in = X"84") then
		sig_out <= X"56";
	elsif (sig_in = X"85") then
		sig_out <= X"57";
	elsif (sig_in = X"86") then
		sig_out <= X"58";
	elsif (sig_in = X"87") then
		sig_out <= X"59";
	elsif (sig_in = X"88") then
		sig_out <= X"5A";
	elsif (sig_in = X"89") then
		sig_out <= X"5B";
	elsif (sig_in = X"8A") then
		sig_out <= X"5C";
	elsif (sig_in = X"8B") then
		sig_out <= X"5D";
	elsif (sig_in = X"8C") then
		sig_out <= X"5E";
	elsif (sig_in = X"8D") then
		sig_out <= X"5F";
	elsif (sig_in = X"8E") then
		sig_out <= X"60";
	elsif (sig_in = X"8F") then
		sig_out <= X"60";
	elsif (sig_in = X"90") then
		sig_out <= X"61";
	elsif (sig_in = X"91") then
		sig_out <= X"62";
	elsif (sig_in = X"92") then
		sig_out <= X"64";
	elsif (sig_in = X"93") then
		sig_out <= X"65";
	elsif (sig_in = X"94") then
		sig_out <= X"66";
	elsif (sig_in = X"95") then
		sig_out <= X"67";
	elsif (sig_in = X"96") then
		sig_out <= X"68";
	elsif (sig_in = X"97") then
		sig_out <= X"69";
	elsif (sig_in = X"98") then
		sig_out <= X"6A";
	elsif (sig_in = X"99") then
		sig_out <= X"6B";
	elsif (sig_in = X"9A") then
		sig_out <= X"6C";
	elsif (sig_in = X"9B") then
		sig_out <= X"6D";
	elsif (sig_in = X"9C") then
		sig_out <= X"6E";
	elsif (sig_in = X"9D") then
		sig_out <= X"6F";
	elsif (sig_in = X"9E") then
		sig_out <= X"70";
	elsif (sig_in = X"9F") then
		sig_out <= X"71";
	elsif (sig_in = X"A0") then
		sig_out <= X"72";
	elsif (sig_in = X"A1") then
		sig_out <= X"73";
	elsif (sig_in = X"A2") then
		sig_out <= X"75";
	elsif (sig_in = X"A3") then
		sig_out <= X"76";
	elsif (sig_in = X"A4") then
		sig_out <= X"77";
	elsif (sig_in = X"A5") then
		sig_out <= X"78";
	elsif (sig_in = X"A6") then
		sig_out <= X"79";
	elsif (sig_in = X"A7") then
		sig_out <= X"7A";
	elsif (sig_in = X"A8") then
		sig_out <= X"7B";
	elsif (sig_in = X"A9") then
		sig_out <= X"7D";
	elsif (sig_in = X"AA") then
		sig_out <= X"7E";
	elsif (sig_in = X"AB") then
		sig_out <= X"7F";
	elsif (sig_in = X"AC") then
		sig_out <= X"80";
	elsif (sig_in = X"AD") then
		sig_out <= X"81";
	elsif (sig_in = X"AE") then
		sig_out <= X"82";
	elsif (sig_in = X"AF") then
		sig_out <= X"84";
	elsif (sig_in = X"B0") then
		sig_out <= X"85";
	elsif (sig_in = X"B1") then
		sig_out <= X"86";
	elsif (sig_in = X"B2") then
		sig_out <= X"87";
	elsif (sig_in = X"B3") then
		sig_out <= X"89";
	elsif (sig_in = X"B4") then
		sig_out <= X"8A";
	elsif (sig_in = X"B5") then
		sig_out <= X"8B";
	elsif (sig_in = X"B6") then
		sig_out <= X"8C";
	elsif (sig_in = X"B7") then
		sig_out <= X"8E";
	elsif (sig_in = X"B8") then
		sig_out <= X"8F";
	elsif (sig_in = X"B9") then
		sig_out <= X"90";
	elsif (sig_in = X"BA") then
		sig_out <= X"91";
	elsif (sig_in = X"BB") then
		sig_out <= X"93";
	elsif (sig_in = X"BC") then
		sig_out <= X"94";
	elsif (sig_in = X"BD") then
		sig_out <= X"95";
	elsif (sig_in = X"BE") then
		sig_out <= X"97";
	elsif (sig_in = X"BF") then
		sig_out <= X"98";
	elsif (sig_in = X"C0") then
		sig_out <= X"99";
	elsif (sig_in = X"C1") then
		sig_out <= X"9B";
	elsif (sig_in = X"C2") then
		sig_out <= X"9C";
	elsif (sig_in = X"C3") then
		sig_out <= X"9D";
	elsif (sig_in = X"C4") then
		sig_out <= X"9F";
	elsif (sig_in = X"C5") then
		sig_out <= X"A0";
	elsif (sig_in = X"C6") then
		sig_out <= X"A2";
	elsif (sig_in = X"C7") then
		sig_out <= X"A3";
	elsif (sig_in = X"C8") then
		sig_out <= X"A4";
	elsif (sig_in = X"C9") then
		sig_out <= X"A6";
	elsif (sig_in = X"CA") then
		sig_out <= X"A7";
	elsif (sig_in = X"CB") then
		sig_out <= X"A9";
	elsif (sig_in = X"CC") then
		sig_out <= X"AA";
	elsif (sig_in = X"CD") then
		sig_out <= X"AB";
	elsif (sig_in = X"CE") then
		sig_out <= X"AD";
	elsif (sig_in = X"CF") then
		sig_out <= X"AE";
	elsif (sig_in = X"D0") then
		sig_out <= X"B0";
	elsif (sig_in = X"D1") then
		sig_out <= X"B1";
	elsif (sig_in = X"D2") then
		sig_out <= X"B3";
	elsif (sig_in = X"D3") then
		sig_out <= X"B4";
	elsif (sig_in = X"D4") then
		sig_out <= X"B6";
	elsif (sig_in = X"D5") then
		sig_out <= X"B7";
	elsif (sig_in = X"D6") then
		sig_out <= X"B9";
	elsif (sig_in = X"D7") then
		sig_out <= X"BA";
	elsif (sig_in = X"D8") then
		sig_out <= X"BC";
	elsif (sig_in = X"D9") then
		sig_out <= X"BD";
	elsif (sig_in = X"DA") then
		sig_out <= X"BF";
	elsif (sig_in = X"DB") then
		sig_out <= X"C1";
	elsif (sig_in = X"DC") then
		sig_out <= X"C2";
	elsif (sig_in = X"DD") then
		sig_out <= X"C4";
	elsif (sig_in = X"DE") then
		sig_out <= X"C5";
	elsif (sig_in = X"DF") then
		sig_out <= X"C7";
	elsif (sig_in = X"E0") then
		sig_out <= X"C8";
	elsif (sig_in = X"E1") then
		sig_out <= X"CA";
	elsif (sig_in = X"E2") then
		sig_out <= X"CC";
	elsif (sig_in = X"E3") then
		sig_out <= X"CD";
	elsif (sig_in = X"E4") then
		sig_out <= X"CF";
	elsif (sig_in = X"E5") then
		sig_out <= X"D1";
	elsif (sig_in = X"E6") then
		sig_out <= X"D2";
	elsif (sig_in = X"E7") then
		sig_out <= X"D4";
	elsif (sig_in = X"E8") then
		sig_out <= X"D6";
	elsif (sig_in = X"E9") then
		sig_out <= X"D7";
	elsif (sig_in = X"EA") then
		sig_out <= X"D9";
	elsif (sig_in = X"EB") then
		sig_out <= X"DB";
	elsif (sig_in = X"EC") then
		sig_out <= X"DC";
	elsif (sig_in = X"ED") then
		sig_out <= X"DE";
	elsif (sig_in = X"EE") then
		sig_out <= X"E0";
	elsif (sig_in = X"EF") then
		sig_out <= X"E2";
	elsif (sig_in = X"F0") then
		sig_out <= X"E3";
	elsif (sig_in = X"F1") then
		sig_out <= X"E5";
	elsif (sig_in = X"F2") then
		sig_out <= X"E7";
	elsif (sig_in = X"F3") then
		sig_out <= X"E9";
	elsif (sig_in = X"F4") then
		sig_out <= X"EA";
	elsif (sig_in = X"F5") then
		sig_out <= X"EC";
	elsif (sig_in = X"F6") then
		sig_out <= X"EE";
	elsif (sig_in = X"F7") then
		sig_out <= X"F0";
	elsif (sig_in = X"F8") then
		sig_out <= X"F2";
	elsif (sig_in = X"F9") then
		sig_out <= X"F4";
	elsif (sig_in = X"FA") then
		sig_out <= X"F5";
	elsif (sig_in = X"FB") then
		sig_out <= X"F7";
	elsif (sig_in = X"FC") then
		sig_out <= X"F9";
	elsif (sig_in = X"FD") then
		sig_out <= X"FB";
	elsif (sig_in = X"FE") then
		sig_out <= X"FD";
	else
		sig_out <= X"FF";
	end if;
	end process;
end architecture;
